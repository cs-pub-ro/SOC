`timescale 1ns / 1ps
module task3(
    output wire o_w_out,
    input wire[1:0] i_w_sel,
    input wire i_w_in1,
    input wire i_w_in2,
    input wire i_w_clk,
    input wire i_w_reset,
    input wire[4:0] i_w_prescaler
);
    
endmodule

module ex1(
    output	out,
    input	in
    );

    not(out, in);
	
endmodule
